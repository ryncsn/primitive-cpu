module Step_Timer_CLR(t0,t1,t2,t3,t4,t5,t6,t7,t8,t9,t10,t11,T_0,T_1,CLK);
input T_0,T_1,CLK;
output t0,t1,t2,t3,t4,t5,t6,t7,t8,t9,t10,t11;
reg t0=1,t1=0,t2=0,t3=0,t4=0,t5=0,t6=0,t7=0,t8=0,t9=0,t10=0,t11=0;
always@(negedge CLK)
begin
if(T_0==1)
{t11,t10,t9,t8,t7,t6,t5,t4,t3,t2,t1,t0}=12'b0000000000000001;
else
if(T_1==1)
begin
case({t11,t10,t9,t8,t7,t6,t5,t4,t3,t2,t1,t0})
12'b000000000001:{t11,t10,t9,t8,t7,t6,t5,t4,t3,t2,t1,t0}=12'b000000000010;
12'b000000000010:{t11,t10,t9,t8,t7,t6,t5,t4,t3,t2,t1,t0}=12'b000000000100;
12'b000000000100:{t11,t10,t9,t8,t7,t6,t5,t4,t3,t2,t1,t0}=12'b000000001000;
12'b000000001000:{t11,t10,t9,t8,t7,t6,t5,t4,t3,t2,t1,t0}=12'b000000010000;
12'b000000010000:{t11,t10,t9,t8,t7,t6,t5,t4,t3,t2,t1,t0}=12'b000000100000;
12'b000000100000:{t11,t10,t9,t8,t7,t6,t5,t4,t3,t2,t1,t0}=12'b000001000000;
12'b000001000000:{t11,t10,t9,t8,t7,t6,t5,t4,t3,t2,t1,t0}=12'b000010000000;
12'b000010000000:{t11,t10,t9,t8,t7,t6,t5,t4,t3,t2,t1,t0}=12'b000100000000;
12'b000100000000:{t11,t10,t9,t8,t7,t6,t5,t4,t3,t2,t1,t0}=12'b001000000000;
12'b001000000000:{t11,t10,t9,t8,t7,t6,t5,t4,t3,t2,t1,t0}=12'b010000000000;
12'b010000000000:{t11,t10,t9,t8,t7,t6,t5,t4,t3,t2,t1,t0}=12'b100000000000;
12'b100000000000:{t11,t10,t9,t8,t7,t6,t5,t4,t3,t2,t1,t0}=12'b000000000001;
default:{t11,t10,t9,t8,t7,t6,t5,t4,t3,t2,t1,t0}=12'b000000000001;
endcase
end
end
endmodule 